library verilog;
use verilog.vl_types.all;
entity test_sum8r is
end test_sum8r;
