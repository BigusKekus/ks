library verilog;
use verilog.vl_types.all;
entity tb_mux4to1_8bit is
end tb_mux4to1_8bit;
